class router_source_sequencer extends uvm_sequencer #(source_xtn);

// Factory registration using `uvm_component_utils
	`uvm_component_utils(router_source_sequencer)

//------------------------------------------
// METHODS
//------------------------------------------

// Standard UVM Methods:
	extern function new(string name = "router_source_sequencer",uvm_component parent);
	endclass
//-----------------  constructor new method  -------------------//
	function router_source_sequencer::new(string name="router_source_sequencer",uvm_component parent);
		super.new(name,parent);
	endfunction



